`timescale 1ns / 1ps

module Delay_op(
    input wire clk,
    input wire rst,
    input wire [10:0] hcount,
    input wire [9:0] vcount,
    input wire hblnk,
    input wire vblnk,
    input wire hsync,
    input wire vsync,
    input wire [11:0] xpos,
    input wire [11:0] ypos,
    
    output reg [10:0] hcount_out,
    output reg [9:0] vcount_out,
    output reg hblnk_out,
    output reg vblnk_out,
    output reg hsync_out,
    output reg vsync_out,
    output reg [11:0] xpos_out,
    output reg [11:0] ypos_out  
    );  
    
    always@(posedge clk)
        if(rst) begin
            hsync_out <= 0;
            vsync_out <= 0;
            hblnk_out <= 0;
            vblnk_out <= 0;
            hcount_out <= 0;
            vcount_out <= 0;
            xpos_out <= xpos;
            ypos_out <= ypos;
        end
        else begin
            hsync_out <= hsync;
            vsync_out <= vsync;
            hblnk_out <= hblnk;
            vblnk_out <= vblnk;
            hcount_out <= hcount;
            vcount_out <= vcount;

            xpos_out <= xpos;
            ypos_out <= ypos;
        end
endmodule
